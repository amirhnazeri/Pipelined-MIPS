`timescale 1ns/1ns

module TestBench();
   reg clk = 0, rst = 0;
   reg[31:0] instMemory[0:65535];
   reg[31:0] regMem[0:31];
   Main uut(clk, rst, instMemory, regMem);

   always #23 clk = ~clk;
   integer i;
   initial begin
      regMem[0] = 32'b00000000000000000000000000000000;
      regMem[1] = 32'b00000000000000000000000000000001;
      regMem[2] = 32'b00000000000000000000000000000010;
      regMem[3] = 32'b00000000000000000000000000000011;
      regMem[4] = 32'b00000000000000000000000000000100;
      regMem[5] = 32'b00000000000000000000000000000101;
      regMem[6] = 32'b00000000000000000000000000000110;
      regMem[7] = 32'b00000000000000000000000000000111;
      regMem[8] = 32'b00000000000000000000000000001000; 
      regMem[9] = 32'b00000000000000000000000000001001; 
      regMem[10] = 32'b00000000000000000000000000001010;
      regMem[11] = 32'b00000000000000000000000000000001;
      regMem[12] = 32'b00000000000000000000000000000010;
      regMem[13] = 32'b00000000000000000000000000000011;
      regMem[14] = 32'b00000000000000000000000000000100;
      regMem[15] = 32'b00000000000000000000000000000101;
      regMem[16] = 32'b00000000000000000000000000000110;
      regMem[17] = 32'b00000000000000000000000000000111;
      regMem[18] = 32'b00000000000000000000000000001000; 
      regMem[19] = 32'b00000000000000000000000000001001; 
      regMem[20] = 32'b00000000000000000000000000001010;
      regMem[21] = 32'b00000000000000000000000000000001;
      regMem[22] = 32'b00000000000000000000000000000001;
      regMem[23] = 32'b00000000000000000000000000000000;
      regMem[24] = 32'b00000000000000000000000000000000;
      regMem[25] = 32'b00000000000000000000000000000000;
      regMem[26] = 32'b00000000000000000000000000000000;
      regMem[27] = 32'b00000000000000000000000000000000;
      regMem[28] = 32'b00000000000000000000000000000000;
      regMem[29] = 32'b00000000000000000000000000000000;
      regMem[30] = 32'b00000000000000000000000000000000;
      regMem[31] = 32'b00000000000000000000000000000000;

      instMemory[0] = 32'b10101100000000010000001111101000; // mem[R0 + 1000] = R1
      instMemory[1] = 32'b10101100000000010000011111010000; // mem[R0 + 2000] = R1
      instMemory[2] = 32'b10001100000101010000001111101000; // R21 = mem[R0 + 1000]
      instMemory[3] = 32'b10001100000101100000011111010000; // R22 = mem[R0 + 2000]
      instMemory[4] = 32'b00000010101101101011100000100000; // R23 = R21 + R22
      
      instMemory[6] = 32'b10101100000000100000001111101001; // mem[R0 + 1001] = R2
      instMemory[7] = 32'b10101100000000100000011111010001; // mem[R0 + 2001] = R2
      instMemory[8] = 32'b10001100000101010000001111101001; // R21 = mem[R0 + 1001]
      instMemory[9] = 32'b10001100000101100000011111010001; // R22 = mem[R0 + 2001]
      instMemory[10] = 32'b00000010101101101011100000100000; // R23 = R21 + R22
      instMemory[11] = 32'b10101100000101110000101110111000; // mem[R0 + 3000] = R23
      
      instMemory[12] = 32'b10101100000000110000001111101010; // mem[R0 + 1002] = R3
      instMemory[13] = 32'b10101100000000110000011111010010; // mem[R0 + 2002] = R3
      instMemory[14] = 32'b10001100000101010000001111101010; // R21 = mem[R0 + 1002]
      instMemory[15] = 32'b10001100000101100000011111010010; // R22 = mem[R0 + 2002]
      instMemory[16] = 32'b00000010101101101011100000100000; // R23 = R21 + R22
      instMemory[17] = 32'b10101100000101110000101110111001; // mem[R0 + 3001] = R23
      
      instMemory[18] = 32'b10101100000001000000001111101011; // mem[R0 + 1003] = R4
      instMemory[19] = 32'b10101100000001000000011111010011; // mem[R0 + 2003] = R4
      instMemory[20] = 32'b10001100000101010000001111101011; // R21 = mem[R0 + 1003]
      instMemory[21] = 32'b10001100000101100000011111010011; // R22 = mem[R0 + 2003]
      instMemory[22] = 32'b00000010101101101011100000100000; // R23 = R21 + R22
      instMemory[23] = 32'b10101100000101110000101110111010; // mem[R0 + 3002] = R23
      
      instMemory[24] = 32'b10101100000001010000001111101100; // mem[R0 + 1004] = R5
      instMemory[25] = 32'b10101100000001010000011111010100; // mem[R0 + 2004] = R5
      instMemory[26] = 32'b10001100000101010000001111101100; // R21 = mem[R0 + 1004]
      instMemory[27] = 32'b10001100000101100000011111010100; // R22 = mem[R0 + 2004]
      instMemory[28] = 32'b00000010101101101011100000100000; // R23 = R21 + R22
      instMemory[29] = 32'b10101100000101110000101110111011; // mem[R0 + 3003] = R23
      
      instMemory[30] = 32'b10101100000001100000001111101101; // mem[R0 + 1005] = R6
      instMemory[31] = 32'b10101100000001100000011111010101; // mem[R0 + 2005] = R6
      instMemory[32] = 32'b10001100000101010000001111101101; // R21 = mem[R0 + 1005]
      instMemory[33] = 32'b10001100000101100000011111010101; // R22 = mem[R0 + 2005]
      instMemory[34] = 32'b00000010101101101011100000100000; // R23 = R21 + R22
      instMemory[35] = 32'b10101100000101110000101110111100; // mem[R0 + 3004] = R23
      
      instMemory[36] = 32'b10101100000001110000001111101110; // mem[R0 + 1006] = R7
      instMemory[37] = 32'b10101100000001110000011111010110; // mem[R0 + 2006] = R7
      instMemory[38] = 32'b10001100000101010000001111101110; // R21 = mem[R0 + 1006]
      instMemory[39] = 32'b10001100000101100000011111010110; // R22 = mem[R0 + 2006]
      instMemory[40] = 32'b00000010101101101011100000100000; // R23 = R21 + R22
      instMemory[41] = 32'b10101100000101110000101110111101; // mem[R0 + 3005] = R23
      
      instMemory[42] = 32'b10101100000010000000001111101111; // mem[R0 + 1007] = R8
      instMemory[43] = 32'b10101100000010000000011111010111; // mem[R0 + 2007] = R8
      instMemory[44] = 32'b10001100000101010000001111101111; // R21 = mem[R0 + 1007]
      instMemory[45] = 32'b10001100000101100000011111010111; // R22 = mem[R0 + 2007]
      instMemory[46] = 32'b00000010101101101011100000100000; // R23 = R21 + R22
      instMemory[47] = 32'b10101100000101110000101110111110; // mem[R0 + 3006] = R23
      
      instMemory[48] = 32'b10101100000010010000001111110000; // mem[R0 + 1008] = R9
      instMemory[49] = 32'b10101100000010010000011111011000; // mem[R0 + 2008] = R9
      instMemory[50] = 32'b10001100000101010000001111110000; // R21 = mem[R0 + 1008]
      instMemory[51] = 32'b10001100000101100000011111011000; // R22 = mem[R0 + 2008]
      instMemory[52] = 32'b00000010101101101011100000100000; // R23 = R21 + R22
      instMemory[53] = 32'b10101100000101110000101110111111; // mem[R0 + 3007] = R23
      
      instMemory[54] = 32'b10101100000010100000001111110001; // mem[R0 + 1009] = R10
      instMemory[55] = 32'b10101100000010100000011111011001; // mem[R0 + 2009] = R10
      instMemory[56] = 32'b10001100000101010000001111110001; // R21 = mem[R0 + 1009]
      instMemory[57] = 32'b10001100000101100000011111011001; // R22 = mem[R0 + 2009]
      instMemory[58] = 32'b00000010101101101011100000100000; // R23 = R21 + R22
      instMemory[59] = 32'b10101100000101110000101111000000; // mem[R0 + 3008] = R23
      
      instMemory[60] = 32'b10101100000010100000001111110001; // mem[R0 + 1009] = R10
      instMemory[61] = 32'b10101100000010100000011111011001; // mem[R0 + 2009] = R10
      instMemory[62] = 32'b10001100000101010000001111110001; // R21 = mem[R0 + 1009]
      instMemory[63] = 32'b10001100000101100000011111011001; // R22 = mem[R0 + 2009]
      instMemory[64] = 32'b00000010101101101011100000100000; // R23 = R21 + R22
      instMemory[65] = 32'b10101100000101110000101111000001; // mem[R0 + 3009] = R23
      
      for(i=66  ; i < 65536; i=i+1) instMemory[i] = 32'b00000000000000000000000000000000;

      rst = 1'b1;
      #85 rst = 1'b0;
      #5850 $stop();
   end
endmodule





